----------------------------------------------------------------------------------
-- Company: 
-- Engineer: Lucia Brown
-- 
-- Create Date: 11/20/2023 08:19:26 PM
-- Design Name: 
-- Module Name: CPU_ControlMemory_22336688 - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
entity CPU_ControlMemory_22336688 is
Port (
Address : in std_logic_vector(16 downto 0);
FL : out std_logic;
FS : out std_logic_vector (4 downto 0);
IL : out std_logic;
MB : out std_logic;
MC : out std_logic;
MD : out std_logic;
MM : out std_logic;
MS : out std_logic_vector (2 downto 0);
MW : out std_logic;
NA : out std_logic_vector (16 downto 0);
PI : out std_logic;
PL : out std_logic;
RC : out std_logic;
RN : out std_logic;
RW : out std_logic;
RV : out std_logic;
RZ : out std_logic;
TA : out std_logic_vector (3 downto 0);
TB : out std_logic_vector (3 downto 0);
TD : out std_logic_vector (3 downto 0)
 );
end CPU_ControlMemory_22336688;

architecture Behavioral of CPU_ControlMemory_22336688 is
-- we u s e t h e l e a s t s i g n i f i c a n t 7 b i t o f t h e Add r e s s - a r r a y ( 0 t o 1 2 7 )
 type ROM_array is array ( 0 to 127 ) of STD_LOGIC_VECTOR ( 50 downto 0 ) ;

 signal ROM : ROM_array := (

 --|5 0 3 4|3 3 3 1 | 3 0 | 2 9| 2 8| 2 7|2 6 2 3|2 2 1 9|1 8 1 5| 1 4|1 3 0 9| 0 8| 0 7| 0 6| 0 5| 0 4| 0 3| 0 2| 0 1| 0 0| C o n t r o l Memory
 --| Next Add r e s s | MS |MC| IL | PI | PL | TD | TA | TB | MB| FS | MD| RW| MM| MW| RV| RC| RN| RZ| FL | Add r e s s
"00000000001011000" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '0' & '1' & '0' & '1' & '1' & '0' & '0' & '0', -- 00 /88
"00000000001011001" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '0' & '1' & '0' & '1' & '1' & '0' & '0' & '1', -- 01 /89
"00000000001011010" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '0' & '1' & '0' & '1' & '1' & '0' & '1' & '0', -- 02 /90
"00000000001011011" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '0' & '1' & '0' & '1' & '1' & '0' & '1' & '1', -- 03 /91
"00000000001011100" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '0' & '1' & '0' & '1' & '1' & '1' & '0' & '0', -- 04 /92
"00000000001011101" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '0' & '1' & '0' & '1' & '1' & '1' & '0' & '1', -- 05 /93
"00000000001011110" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '0' & '1' & '0' & '1' & '1' & '1' & '1' & '0', -- 06 /94
"00000000001011111" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '0' & '1' & '0' & '1' & '1' & '1' & '1' & '1', -- 07 /95
"00000000001100000" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '0' & '1' & '1' & '0' & '0' & '0' & '0' & '0', -- 08 /96
"00000000001100001" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '0' & '1' & '1' & '0' & '0' & '0' & '0' & '1', -- 09 /97
"00000000001100010" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '0' & '1' & '1' & '0' & '0' & '0' & '1' & '0', -- 0A /98
"00000000001100011" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '0' & '1' & '1' & '0' & '0' & '0' & '1' & '1', -- 0B /99
"00000000001100100" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '0' & '1' & '1' & '0' & '0' & '1' & '0' & '0', -- 0C /100
"00000000001100101" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '0' & '1' & '1' & '0' & '0' & '1' & '0' & '1', -- 0D /101
"00000000001100110" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '0' & '1' & '1' & '0' & '0' & '1' & '1' & '0', -- 0E /102
"00000000001100111" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '0' & '1' & '1' & '0' & '0' & '1' & '1' & '1', -- 0F /103


"00000000001101000" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '0' & '1' & '1' & '0' & '1' & '0' & '0' & '0', -- 10 /104
"00000000001101001" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '0' & '1' & '1' & '0' & '1' & '0' & '0' & '1', -- 11 /105
"00000000001101010" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '0' & '1' & '1' & '0' & '1' & '0' & '1' & '0', -- 12 /106
"00000000001101011" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '0' & '1' & '1' & '0' & '1' & '0' & '1' & '1', -- 13 /107
"00000000001101100" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '0' & '1' & '1' & '0' & '1' & '1' & '0' & '0', -- 14 /108
"00000000001101101" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '0' & '1' & '1' & '0' & '1' & '1' & '0' & '1', -- 15 /109
"00000000001101110" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '0' & '1' & '1' & '0' & '1' & '1' & '1' & '0', -- 16 /110
"00000000001101111" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '0' & '1' & '1' & '0' & '1' & '1' & '1' & '1', -- 17 /111
"00000000001110000" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '0' & '1' & '1' & '1' & '0' & '0' & '0' & '0', -- 18 /112
"00000000001110001" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '0' & '1' & '1' & '1' & '0' & '0' & '0' & '1', -- 19 /113
"00000000001110010" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '0' & '1' & '1' & '1' & '0' & '0' & '1' & '0', -- 1A /114
"00000000001110011" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '0' & '1' & '1' & '1' & '0' & '0' & '1' & '1', -- 1B /115
"00000000001110100" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '0' & '1' & '1' & '1' & '0' & '1' & '0' & '0', -- 1C /116
"00000000001110101" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '0' & '1' & '1' & '1' & '0' & '1' & '0' & '1', -- 1D /117
"00000000001110110" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '0' & '1' & '1' & '1' & '0' & '1' & '1' & '0', -- 1E /118
"00000000001110111" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '0' & '1' & '1' & '1' & '0' & '1' & '1' & '1', -- 1F /119


 --|5 0 3 4|3 3 3 1 | 3 0 | 2 9| 2 8| 2 7|2 6 2 3|2 2 1 9|1 8 1 5| 1 4|1 3 0 9| 0 8| 0 7| 0 6| 0 5| 0 4| 0 3| 0 2| 0 1| 0 0| C o n t r o l Memory
 --| Next Add r e s s | MS |MC| IL | PI | PL | TD | TA | TB | MB| FS | MD| RW| MM| MW| RV| RC| RN| RZ| FL | Add r e s s
"00000000001111000" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '0' & '1' & '1' & '1' & '1' & '0' & '0' & '0', -- 20/120
"00000000001111001" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '0' & '1' & '1' & '1' & '1' & '0' & '0' & '1', -- 21/121
"00000000001111010" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '0' & '1' & '1' & '1' & '1' & '0' & '1' & '0', -- 22/122
"00000000001111011" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '0' & '1' & '1' & '1' & '1' & '0' & '1' & '1', -- 23/123
"00000000001111100" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '0' & '1' & '1' & '1' & '1' & '1' & '0' & '0', -- 24/124
"00000000001111101" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '0' & '1' & '1' & '1' & '1' & '1' & '0' & '1', -- 25/125
"00000000001111110" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '0' & '1' & '1' & '1' & '1' & '1' & '1' & '0', -- 26/126
"00000000001111111" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '0' & '1' & '1' & '1' & '1' & '1' & '1' & '1', -- 27/127
"00000000010000000" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '1' & '0' & '0' & '0' & '0' & '0' & '0' & '0', -- 28/128
"00000000010000001" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '1' & '0' & '0' & '0' & '0' & '0' & '0' & '1', -- 29/129
"00000000010000010" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '1' & '0' & '0' & '0' & '0' & '0' & '1' & '0', -- 2A/130
"00000000010000011" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '1' & '0' & '0' & '0' & '0' & '0' & '1' & '1', -- 2B/131
"00000000010000100" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '1' & '0' & '0' & '0' & '0' & '1' & '0' & '0', -- 2C/132
"00000000010000101" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '1' & '0' & '0' & '0' & '0' & '1' & '0' & '1', -- 2D/133
"00000000010000110" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '1' & '0' & '0' & '0' & '0' & '1' & '1' & '0', -- 2E/134
"00000000010000111" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '1' & '0' & '0' & '0' & '0' & '1' & '1' & '1',  -- 2F/135

--|5 0 3 4|3 3 3 1 | 3 0 | 2 9| 2 8| 2 7|2 6 2 3|2 2 1 9|1 8 1 5| 1 4|1 3 0 9| 0 8| 0 7| 0 6| 0 5| 0 4| 0 3| 0 2| 0 1| 0 0| C o n t r o l Memory
--| Next Add r e s s | MS |MC| IL | PI | PL | TD | TA | TB | MB| FS | MD| RW| MM| MW| RV| RC| RN| RZ| FL | Add r e s s
"00000000010001000" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '1' & '0' & '0' & '0' & '1' & '0' & '0' & '0', -- 30/136
"00000000010001001" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '1' & '0' & '0' & '0' & '1' & '0' & '0' & '1', -- 31/137
"00000000010001010" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '1' & '0' & '0' & '0' & '1' & '0' & '1' & '0', -- 32/138
"00000000010001011" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '1' & '0' & '0' & '0' & '1' & '0' & '1' & '1', -- 33/139
"00000000010001100" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '1' & '0' & '0' & '0' & '1' & '1' & '0' & '0', -- 34/140
"00000000010001101" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '1' & '0' & '0' & '0' & '1' & '1' & '0' & '1', -- 35/141
"00000000010001110" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '1' & '0' & '0' & '0' & '1' & '1' & '1' & '0', -- 36/142
"00000000010001111" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '1' & '0' & '0' & '0' & '1' & '1' & '1' & '1', -- 37/143
"00000000010010000" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '1' & '0' & '0' & '1' & '0' & '0' & '0' & '0', -- 38/144
"00000000010010001" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '1' & '0' & '0' & '1' & '0' & '0' & '0' & '1', -- 39/145
"00000000010010010" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '1' & '0' & '0' & '1' & '0' & '0' & '1' & '0', -- 3A/146
"00000000010010011" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '1' & '0' & '0' & '1' & '0' & '0' & '1' & '1', -- 3B/147
"00000000010010100" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '1' & '0' & '0' & '1' & '0' & '1' & '0' & '0', -- 3C/148
"00000000010010101" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '1' & '0' & '0' & '1' & '0' & '1' & '0' & '1', -- 3D/149
"00000000010010110" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '1' & '0' & '0' & '1' & '0' & '1' & '1' & '0', -- 3E/150
"00000000010010111" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '1' & '0' & '0' & '1' & '0' & '1' & '1' & '1',  -- 3F/151




 --|5 0 3 4|3 3 3 1 | 3 0 | 2 9| 2 8| 2 7|2 6 2 3|2 2 1 9|1 8 1 5| 1 4|1 3 0 9| 0 8| 0 7| 0 6| 0 5| 0 4| 0 3| 0 2| 0 1| 0 0| C o n t r o l Memory
 --| Next Add r e s s | MS |MC| IL | PI | PL | TD | TA | TB | MB| FS | MD| RW| MM| MW| RV| RC| RN| RZ| FL | Add r e s s
"00000000010011000" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '1' & '0' & '0' & '1' & '1' & '0' & '0' & '0', -- 40/152
"00000000010011001" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '1' & '0' & '0' & '1' & '1' & '0' & '0' & '1', -- 41/153
"00000000010011010" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '1' & '0' & '0' & '1' & '1' & '0' & '1' & '0', -- 42/154
"00000000010011011" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '1' & '0' & '0' & '1' & '1' & '0' & '1' & '1', -- 43/155
"00000000010011100" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '1' & '0' & '0' & '1' & '1' & '1' & '0' & '0', -- 44/156
"00000000010011101" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '1' & '0' & '0' & '1' & '1' & '1' & '0' & '1', -- 45/157
"00000000010011110" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '1' & '0' & '0' & '1' & '1' & '1' & '1' & '0', -- 46/158
"00000000010011111" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '1' & '0' & '0' & '1' & '1' & '1' & '1' & '1', -- 47/159
"00000000010100000" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '1' & '0' & '1' & '0' & '0' & '0' & '0' & '0', -- 48/160
"00000000010100001" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '1' & '0' & '1' & '0' & '0' & '0' & '0' & '1', -- 49/161
"00000000010100010" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '1' & '0' & '1' & '0' & '0' & '0' & '1' & '0', -- 4A/162
"00000000010100011" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '1' & '0' & '1' & '0' & '0' & '0' & '1' & '1', -- 4B/163
"00000000010100100" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '1' & '0' & '1' & '0' & '0' & '1' & '0' & '0', -- 4C/164
"00000000010100101" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '1' & '0' & '1' & '0' & '0' & '1' & '0' & '1', -- 4D/165
"00000000010100110" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '1' & '0' & '1' & '0' & '0' & '1' & '1' & '0', -- 4E/166
"00000000010100111" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '1' & '0' & '1' & '0' & '0' & '1' & '1' & '1',  -- 4F/167



 --|5 0 3 4|3 3 3 1 | 3 0 | 2 9| 2 8| 2 7|2 6 2 3|2 2 1 9|1 8 1 5| 1 4|1 3 0 9| 0 8| 0 7| 0 6| 0 5| 0 4| 0 3| 0 2| 0 1| 0 0| C o n t r o l Memory
 --| Next Add r e s s | MS |MC| IL | PI | PL | TD | TA | TB | MB| FS | MD| RW| MM| MW| RV| RC| RN| RZ| FL | Add r e s s
"00000000010101000" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '1' & '0' & '1' & '0' & '1' & '0' & '0' & '0', -- 50/168
"00000000010101001" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '1' & '0' & '1' & '0' & '1' & '0' & '0' & '1', -- 51/169
"00000000010101010" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '1' & '0' & '1' & '0' & '1' & '0' & '1' & '0', -- 52/170
"00000000010101011" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '1' & '0' & '1' & '0' & '1' & '0' & '1' & '1', -- 53/171
"00000000010101100" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '1' & '0' & '1' & '0' & '1' & '1' & '0' & '0', -- 54/172
"00000000010101101" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '1' & '0' & '1' & '0' & '1' & '1' & '0' & '1', -- 55/173
"00000000010101110" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '1' & '0' & '1' & '0' & '1' & '1' & '1' & '0', -- 56/174
"00000000010101111" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '1' & '0' & '1' & '0' & '1' & '1' & '1' & '1', -- 57/175
"00000000010110000" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '1' & '0' & '1' & '1' & '0' & '0' & '0' & '0', -- 58/176
"00000000010110001" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '1' & '0' & '1' & '1' & '0' & '0' & '0' & '1', -- 59/177
"00000000010110010" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '1' & '0' & '1' & '1' & '0' & '0' & '1' & '0', -- 5A/178
"00000000010110011" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '1' & '0' & '1' & '1' & '0' & '0' & '1' & '1', -- 5B/179
"00000000010110100" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '1' & '0' & '1' & '1' & '0' & '1' & '0' & '0', -- 5C/180
"00000000010110101" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '1' & '0' & '1' & '1' & '0' & '1' & '0' & '1', -- 5D/181
"00000000010110110" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '1' & '0' & '1' & '1' & '0' & '1' & '1' & '0', -- 5E/182
"00000000010110111" & "000" & '0' & '0' & '0' & '0' & "0000" & "0000" & "0000" & '0' & "00000" & '0' & '1' & '0' & '1' & '1' & '0' & '1' & '1' & '1',  -- 5F/183




 --|5 0 3 4|3 3 3 1 | 3 0 | 2 9| 2 8| 2 7|2 6 2 3|2 2 1 9|1 8 1 5| 1 4|1 3 0 9| 0 8| 0 7| 0 6| 0 5| 0 4| 0 3| 0 2| 0 1| 0 0| C o n t r o l Memory
 --| Next Add r e s s | MS |MC| IL | PI | PL | TD | TA | TB | MB| FS | MD| RW| MM| MW| RV| RC| RN| RZ| FL | Add r e s s
"00000000010111000"&"000" & '0'& '0'& '0'& '0'& "0000"&"0000"&"0000"&'0'&"00000" & '0'& '1'& '0'& '1'& '1'& '1'& '0'& '0'& '0', -- 60/184
"00000000010111001"&"000" & '0'& '0'& '0'& '0'& "0000"&"0000"&"0000"&'0'&"00000" & '0'& '1'& '0'& '1'& '1'& '1'& '0'& '0'& '1', -- 61/185
"00000000010111010"&"000" & '0'& '0'& '0'& '0'& "0000"&"0000"&"0000"&'0'&"00000" & '0'& '1'& '0'& '1'& '1'& '1'& '0'& '1'& '0', -- 62/186
"00000000010111011"&"000" & '0'& '0'& '0'& '0'& "0000"&"0000"&"0000"&'0'&"00000" & '0'& '1'& '0'& '1'& '1'& '1'& '0'& '1'& '1', -- 63/187
"00000000010111100"&"000" & '0'& '0'& '0'& '0'& "0000"&"0000"&"0000"&'0'&"00000" & '0'& '1'& '0'& '1'& '1'& '1'& '1'& '0'& '0', -- 64/188
"00000000010111101"&"000" & '0'& '0'& '0'& '0'& "0000"&"0000"&"0000"&'0'&"00000" & '0'& '1'& '0'& '1'& '1'& '1'& '1'& '0'& '1', -- 65/189
"00000000010111110"&"000" & '0'& '0'& '0'& '0'& "0000"&"0000"&"0000"&'0'&"00000" & '0'& '1'& '0'& '1'& '1'& '1'& '1'& '1'& '0', -- 66/190
"00000000010111111"&"000" & '0'& '0'& '0'& '0'& "0000"&"0000"&"0000"&'0'&"00000" & '0'& '1'& '0'& '1'& '1'& '1'& '1'& '1'& '1', -- 67/191
"00000000011000000"&"000" & '0'& '0'& '0'& '0'& "0000"&"0000"&"0000"&'0'&"00000" & '0'& '1'& '1'& '0'& '0'& '0'& '0'& '0'& '0', -- 68/192
"00000000011000001"&"000" & '0'& '0'& '0'& '0'& "0000"&"0000"&"0000"&'0'&"00000" & '0'& '1'& '1'& '0'& '0'& '0'& '0'& '0'& '1', -- 69/193
"00000000011000010"&"000" & '0'& '0'& '0'& '0'& "0000"&"0000"&"0000"&'0'&"00000" & '0'& '1'& '1'& '0'& '0'& '0'& '0'& '1'& '0', -- 6A/194
"00000000011000011"&"000" & '0'& '0'& '0'& '0'& "0000"&"0000"&"0000"&'0'&"00000" & '0'& '1'& '1'& '0'& '0'& '0'& '0'& '1'& '1', -- 6B/195
"00000000011000100"&"000" & '0'& '0'& '0'& '0'& "0000"&"0000"&"0000"&'0'&"00000" & '0'& '1'& '1'& '0'& '0'& '0'& '1'& '0'& '0', -- 6C/196
"00000000011000101"&"000" & '0'& '0'& '0'& '0'& "0000"&"0000"&"0000"&'0'&"00000" & '0'& '1'& '1'& '0'& '0'& '0'& '1'& '0'& '1', -- 6D/197
"00000000011000110"&"000" & '0'& '0'& '0'& '0'& "0000"&"0000"&"0000"&'0'&"00000" & '0'& '1'& '1'& '0'& '0'& '0'& '1'& '1'& '0', -- 6E/198
"00000000011000111"&"000" & '0'& '0'& '0'& '0'& "0000"&"0000"&"0000"&'0'&"00000" & '0'& '1'& '1'& '0'& '0'& '0'& '1'& '1'& '1', -- 6F/199

 --|5 0 3 4|3 3 3 1 | 3 0 | 2 9| 2 8| 2 7|2 6 2 3|2 2 1 9|1 8 1 5| 1 4|1 3 0 9| 0 8| 0 7| 0 6| 0 5| 0 4| 0 3| 0 2| 0 1| 0 0| C o n t r o l Memory
 --| Next Add r e s s | MS |MC| IL | PI | PL | TD | TA | TB | MB| FS | MD| RW| MM| MW| RV| RC| RN| RZ| FL | Add r e s s
"00000000011001000"&"000" & '0'& '0'& '0'& '0'& "0000"&"0000"&"0000"&'0'&"00000" & '0'& '1'& '1'& '0'& '0'& '1'& '0'& '0'& '0', -- 70/200
"00000000011001001"&"000" & '0'& '0'& '0'& '0'& "0000"&"0000"&"0000"&'0'&"00000" & '0'& '1'& '1'& '0'& '0'& '1'& '0'& '0'& '1', -- 71/201
"00000000011001010"&"000" & '0'& '0'& '0'& '0'& "0000"&"0000"&"0000"&'0'&"00000" & '0'& '1'& '1'& '0'& '0'& '1'& '0'& '1'& '0', -- 72/202
"00000000011001011"&"000" & '0'& '0'& '0'& '0'& "0000"&"0000"&"0000"&'0'&"00000" & '0'& '1'& '1'& '0'& '0'& '1'& '0'& '1'& '1', -- 73/203
"00000000011001100"&"000" & '0'& '0'& '0'& '0'& "0000"&"0000"&"0000"&'0'&"00000" & '0'& '1'& '1'& '0'& '0'& '1'& '1'& '0'& '0', -- 74/204
"00000000011001101"&"000" & '0'& '0'& '0'& '0'& "0000"&"0000"&"0000"&'0'&"00000" & '0'& '1'& '1'& '0'& '0'& '1'& '1'& '0'& '1', -- 75/205
"00000000011001110"&"000" & '0'& '0'& '0'& '0'& "0000"&"0000"&"0000"&'0'&"00000" & '0'& '1'& '1'& '0'& '0'& '1'& '1'& '1'& '0', -- 76/206
"00000000011001111"&"000" & '0'& '0'& '0'& '0'& "0000"&"0000"&"0000"&'0'&"00000" & '0'& '1'& '1'& '0'& '0'& '1'& '1'& '1'& '1', -- 77/207
"00000000011010000"&"000" & '0'& '0'& '0'& '0'& "0000"&"0000"&"0000"&'0'&"00000" & '0'& '1'& '1'& '0'& '1'& '0'& '0'& '0'& '0', -- 78/208
"00000000011010001"&"000" & '0'& '0'& '0'& '0'& "0000"&"0000"&"0000"&'0'&"00000" & '0'& '1'& '1'& '0'& '1'& '0'& '0'& '0'& '1', -- 79/209
"00000000011010010"&"000" & '0'& '0'& '0'& '0'& "0000"&"0000"&"0000"&'0'&"00000" & '0'& '1'& '1'& '0'& '1'& '0'& '0'& '1'& '0', -- 7A/210
"00000000011010011"&"000" & '0'& '0'& '0'& '0'& "0000"&"0000"&"0000"&'0'&"00000" & '0'& '1'& '1'& '0'& '1'& '0'& '0'& '1'& '1', -- 7B/211
"00000000011010100"&"000" & '0'& '0'& '0'& '0'& "0000"&"0000"&"0000"&'0'&"00000" & '0'& '1'& '1'& '0'& '1'& '0'& '1'& '0'& '0', -- 7C/212
"00000000011010101"&"000" & '0'& '0'& '0'& '0'& "0000"&"0000"&"0000"&'0'&"00000" & '0'& '1'& '1'& '0'& '1'& '0'& '1'& '0'& '1', -- 7D/213
"00000000011010110"&"000" & '0'& '0'& '0'& '0'& "0000"&"0000"&"0000"&'0'&"00000" & '0'& '1'& '1'& '0'& '1'& '0'& '1'& '1'& '0', -- 7E/214
"00000000011010111"&"000" & '0'& '0'& '0'& '0'& "0000"&"0000"&"0000"&'0'&"00000" & '0'& '1'& '1'& '0'& '1'& '0'& '1'& '1'& '1' -- 7F/215    

 ) ;

signal content_at_address : STD_LOGIC_VECTOR( 50 downto 0 ) ;
begin
content_at_address<= ROM( to_integer(unsigned(Address(6 downto 0 )))) after 2 ns ;
 NA <= content_at_address ( 50 downto 34 ) ; -- 34-50
 MS <= content_at_address ( 33 downto 31 ) ; -- 31-33
 MC <= content_at_address ( 30 ) ; -- 30
 IL <= content_at_address ( 29 ) ; -- 29
 PI <= content_at_address ( 28 ) ; -- 28
 PL <= content_at_address ( 27 ) ; -- 27
 TD <= content_at_address ( 26 downto 23 ) ; -- 23-26
 TA <= content_at_address ( 22 downto 19 ) ; -- 19-22
 TB <= content_at_address ( 18 downto 15 ) ; -- 15-18
 MB <= content_at_address ( 14 ) ; -- 14
 FS <= content_at_address( 13 downto 9 ) ; -- 09-13
 MD <= content_at_address ( 8 ) ; -- 08
 RW <= content_at_address ( 7 ) ; -- 07
 MM <= content_at_address( 6 ) ; -- 06
 MW <= content_at_address( 5 ) ; -- 05
 RV <= content_at_address ( 4 ) ; -- 04
 RC <= content_at_address( 3 ) ; -- 03
 RN <= content_at_address( 2 ) ; -- 02
 RZ <= content_at_address ( 1 ) ; -- 01
 FL <= content_at_address ( 0 ) ; -- 00


end Behavioral;
